xy
z

abs vgmm
